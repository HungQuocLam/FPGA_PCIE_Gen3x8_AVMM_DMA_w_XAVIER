// top_hw.v

// Generated using ACDS version 19.2 57

`timescale 1 ps / 1 ps
module top_hw (
		input  wire [31:0] hip_ctrl_test_in,                //           hip_ctrl.test_in
		input  wire        hip_ctrl_simu_mode_pipe,         //                   .simu_mode_pipe
		input  wire        hip_pipe_sim_pipe_pclk_in,       //           hip_pipe.sim_pipe_pclk_in
		output wire [1:0]  hip_pipe_sim_pipe_rate,          //                   .sim_pipe_rate
		output wire [4:0]  hip_pipe_sim_ltssmstate,         //                   .sim_ltssmstate
		output wire [2:0]  hip_pipe_eidleinfersel0,         //                   .eidleinfersel0
		output wire [2:0]  hip_pipe_eidleinfersel1,         //                   .eidleinfersel1
		output wire [2:0]  hip_pipe_eidleinfersel2,         //                   .eidleinfersel2
		output wire [2:0]  hip_pipe_eidleinfersel3,         //                   .eidleinfersel3
		output wire [2:0]  hip_pipe_eidleinfersel4,         //                   .eidleinfersel4
		output wire [2:0]  hip_pipe_eidleinfersel5,         //                   .eidleinfersel5
		output wire [2:0]  hip_pipe_eidleinfersel6,         //                   .eidleinfersel6
		output wire [2:0]  hip_pipe_eidleinfersel7,         //                   .eidleinfersel7
		output wire [1:0]  hip_pipe_powerdown0,             //                   .powerdown0
		output wire [1:0]  hip_pipe_powerdown1,             //                   .powerdown1
		output wire [1:0]  hip_pipe_powerdown2,             //                   .powerdown2
		output wire [1:0]  hip_pipe_powerdown3,             //                   .powerdown3
		output wire [1:0]  hip_pipe_powerdown4,             //                   .powerdown4
		output wire [1:0]  hip_pipe_powerdown5,             //                   .powerdown5
		output wire [1:0]  hip_pipe_powerdown6,             //                   .powerdown6
		output wire [1:0]  hip_pipe_powerdown7,             //                   .powerdown7
		output wire        hip_pipe_rxpolarity0,            //                   .rxpolarity0
		output wire        hip_pipe_rxpolarity1,            //                   .rxpolarity1
		output wire        hip_pipe_rxpolarity2,            //                   .rxpolarity2
		output wire        hip_pipe_rxpolarity3,            //                   .rxpolarity3
		output wire        hip_pipe_rxpolarity4,            //                   .rxpolarity4
		output wire        hip_pipe_rxpolarity5,            //                   .rxpolarity5
		output wire        hip_pipe_rxpolarity6,            //                   .rxpolarity6
		output wire        hip_pipe_rxpolarity7,            //                   .rxpolarity7
		output wire        hip_pipe_txcompl0,               //                   .txcompl0
		output wire        hip_pipe_txcompl1,               //                   .txcompl1
		output wire        hip_pipe_txcompl2,               //                   .txcompl2
		output wire        hip_pipe_txcompl3,               //                   .txcompl3
		output wire        hip_pipe_txcompl4,               //                   .txcompl4
		output wire        hip_pipe_txcompl5,               //                   .txcompl5
		output wire        hip_pipe_txcompl6,               //                   .txcompl6
		output wire        hip_pipe_txcompl7,               //                   .txcompl7
		output wire [31:0] hip_pipe_txdata0,                //                   .txdata0
		output wire [31:0] hip_pipe_txdata1,                //                   .txdata1
		output wire [31:0] hip_pipe_txdata2,                //                   .txdata2
		output wire [31:0] hip_pipe_txdata3,                //                   .txdata3
		output wire [31:0] hip_pipe_txdata4,                //                   .txdata4
		output wire [31:0] hip_pipe_txdata5,                //                   .txdata5
		output wire [31:0] hip_pipe_txdata6,                //                   .txdata6
		output wire [31:0] hip_pipe_txdata7,                //                   .txdata7
		output wire [3:0]  hip_pipe_txdatak0,               //                   .txdatak0
		output wire [3:0]  hip_pipe_txdatak1,               //                   .txdatak1
		output wire [3:0]  hip_pipe_txdatak2,               //                   .txdatak2
		output wire [3:0]  hip_pipe_txdatak3,               //                   .txdatak3
		output wire [3:0]  hip_pipe_txdatak4,               //                   .txdatak4
		output wire [3:0]  hip_pipe_txdatak5,               //                   .txdatak5
		output wire [3:0]  hip_pipe_txdatak6,               //                   .txdatak6
		output wire [3:0]  hip_pipe_txdatak7,               //                   .txdatak7
		output wire        hip_pipe_txdetectrx0,            //                   .txdetectrx0
		output wire        hip_pipe_txdetectrx1,            //                   .txdetectrx1
		output wire        hip_pipe_txdetectrx2,            //                   .txdetectrx2
		output wire        hip_pipe_txdetectrx3,            //                   .txdetectrx3
		output wire        hip_pipe_txdetectrx4,            //                   .txdetectrx4
		output wire        hip_pipe_txdetectrx5,            //                   .txdetectrx5
		output wire        hip_pipe_txdetectrx6,            //                   .txdetectrx6
		output wire        hip_pipe_txdetectrx7,            //                   .txdetectrx7
		output wire        hip_pipe_txelecidle0,            //                   .txelecidle0
		output wire        hip_pipe_txelecidle1,            //                   .txelecidle1
		output wire        hip_pipe_txelecidle2,            //                   .txelecidle2
		output wire        hip_pipe_txelecidle3,            //                   .txelecidle3
		output wire        hip_pipe_txelecidle4,            //                   .txelecidle4
		output wire        hip_pipe_txelecidle5,            //                   .txelecidle5
		output wire        hip_pipe_txelecidle6,            //                   .txelecidle6
		output wire        hip_pipe_txelecidle7,            //                   .txelecidle7
		output wire        hip_pipe_txdeemph0,              //                   .txdeemph0
		output wire        hip_pipe_txdeemph1,              //                   .txdeemph1
		output wire        hip_pipe_txdeemph2,              //                   .txdeemph2
		output wire        hip_pipe_txdeemph3,              //                   .txdeemph3
		output wire        hip_pipe_txdeemph4,              //                   .txdeemph4
		output wire        hip_pipe_txdeemph5,              //                   .txdeemph5
		output wire        hip_pipe_txdeemph6,              //                   .txdeemph6
		output wire        hip_pipe_txdeemph7,              //                   .txdeemph7
		output wire [2:0]  hip_pipe_txmargin0,              //                   .txmargin0
		output wire [2:0]  hip_pipe_txmargin1,              //                   .txmargin1
		output wire [2:0]  hip_pipe_txmargin2,              //                   .txmargin2
		output wire [2:0]  hip_pipe_txmargin3,              //                   .txmargin3
		output wire [2:0]  hip_pipe_txmargin4,              //                   .txmargin4
		output wire [2:0]  hip_pipe_txmargin5,              //                   .txmargin5
		output wire [2:0]  hip_pipe_txmargin6,              //                   .txmargin6
		output wire [2:0]  hip_pipe_txmargin7,              //                   .txmargin7
		output wire        hip_pipe_txswing0,               //                   .txswing0
		output wire        hip_pipe_txswing1,               //                   .txswing1
		output wire        hip_pipe_txswing2,               //                   .txswing2
		output wire        hip_pipe_txswing3,               //                   .txswing3
		output wire        hip_pipe_txswing4,               //                   .txswing4
		output wire        hip_pipe_txswing5,               //                   .txswing5
		output wire        hip_pipe_txswing6,               //                   .txswing6
		output wire        hip_pipe_txswing7,               //                   .txswing7
		input  wire        hip_pipe_phystatus0,             //                   .phystatus0
		input  wire        hip_pipe_phystatus1,             //                   .phystatus1
		input  wire        hip_pipe_phystatus2,             //                   .phystatus2
		input  wire        hip_pipe_phystatus3,             //                   .phystatus3
		input  wire        hip_pipe_phystatus4,             //                   .phystatus4
		input  wire        hip_pipe_phystatus5,             //                   .phystatus5
		input  wire        hip_pipe_phystatus6,             //                   .phystatus6
		input  wire        hip_pipe_phystatus7,             //                   .phystatus7
		input  wire [31:0] hip_pipe_rxdata0,                //                   .rxdata0
		input  wire [31:0] hip_pipe_rxdata1,                //                   .rxdata1
		input  wire [31:0] hip_pipe_rxdata2,                //                   .rxdata2
		input  wire [31:0] hip_pipe_rxdata3,                //                   .rxdata3
		input  wire [31:0] hip_pipe_rxdata4,                //                   .rxdata4
		input  wire [31:0] hip_pipe_rxdata5,                //                   .rxdata5
		input  wire [31:0] hip_pipe_rxdata6,                //                   .rxdata6
		input  wire [31:0] hip_pipe_rxdata7,                //                   .rxdata7
		input  wire [3:0]  hip_pipe_rxdatak0,               //                   .rxdatak0
		input  wire [3:0]  hip_pipe_rxdatak1,               //                   .rxdatak1
		input  wire [3:0]  hip_pipe_rxdatak2,               //                   .rxdatak2
		input  wire [3:0]  hip_pipe_rxdatak3,               //                   .rxdatak3
		input  wire [3:0]  hip_pipe_rxdatak4,               //                   .rxdatak4
		input  wire [3:0]  hip_pipe_rxdatak5,               //                   .rxdatak5
		input  wire [3:0]  hip_pipe_rxdatak6,               //                   .rxdatak6
		input  wire [3:0]  hip_pipe_rxdatak7,               //                   .rxdatak7
		input  wire        hip_pipe_rxelecidle0,            //                   .rxelecidle0
		input  wire        hip_pipe_rxelecidle1,            //                   .rxelecidle1
		input  wire        hip_pipe_rxelecidle2,            //                   .rxelecidle2
		input  wire        hip_pipe_rxelecidle3,            //                   .rxelecidle3
		input  wire        hip_pipe_rxelecidle4,            //                   .rxelecidle4
		input  wire        hip_pipe_rxelecidle5,            //                   .rxelecidle5
		input  wire        hip_pipe_rxelecidle6,            //                   .rxelecidle6
		input  wire        hip_pipe_rxelecidle7,            //                   .rxelecidle7
		input  wire [2:0]  hip_pipe_rxstatus0,              //                   .rxstatus0
		input  wire [2:0]  hip_pipe_rxstatus1,              //                   .rxstatus1
		input  wire [2:0]  hip_pipe_rxstatus2,              //                   .rxstatus2
		input  wire [2:0]  hip_pipe_rxstatus3,              //                   .rxstatus3
		input  wire [2:0]  hip_pipe_rxstatus4,              //                   .rxstatus4
		input  wire [2:0]  hip_pipe_rxstatus5,              //                   .rxstatus5
		input  wire [2:0]  hip_pipe_rxstatus6,              //                   .rxstatus6
		input  wire [2:0]  hip_pipe_rxstatus7,              //                   .rxstatus7
		input  wire        hip_pipe_rxvalid0,               //                   .rxvalid0
		input  wire        hip_pipe_rxvalid1,               //                   .rxvalid1
		input  wire        hip_pipe_rxvalid2,               //                   .rxvalid2
		input  wire        hip_pipe_rxvalid3,               //                   .rxvalid3
		input  wire        hip_pipe_rxvalid4,               //                   .rxvalid4
		input  wire        hip_pipe_rxvalid5,               //                   .rxvalid5
		input  wire        hip_pipe_rxvalid6,               //                   .rxvalid6
		input  wire        hip_pipe_rxvalid7,               //                   .rxvalid7
		input  wire        hip_pipe_rxdataskip0,            //                   .rxdataskip0
		input  wire        hip_pipe_rxdataskip1,            //                   .rxdataskip1
		input  wire        hip_pipe_rxdataskip2,            //                   .rxdataskip2
		input  wire        hip_pipe_rxdataskip3,            //                   .rxdataskip3
		input  wire        hip_pipe_rxdataskip4,            //                   .rxdataskip4
		input  wire        hip_pipe_rxdataskip5,            //                   .rxdataskip5
		input  wire        hip_pipe_rxdataskip6,            //                   .rxdataskip6
		input  wire        hip_pipe_rxdataskip7,            //                   .rxdataskip7
		input  wire        hip_pipe_rxblkst0,               //                   .rxblkst0
		input  wire        hip_pipe_rxblkst1,               //                   .rxblkst1
		input  wire        hip_pipe_rxblkst2,               //                   .rxblkst2
		input  wire        hip_pipe_rxblkst3,               //                   .rxblkst3
		input  wire        hip_pipe_rxblkst4,               //                   .rxblkst4
		input  wire        hip_pipe_rxblkst5,               //                   .rxblkst5
		input  wire        hip_pipe_rxblkst6,               //                   .rxblkst6
		input  wire        hip_pipe_rxblkst7,               //                   .rxblkst7
		input  wire [1:0]  hip_pipe_rxsynchd0,              //                   .rxsynchd0
		input  wire [1:0]  hip_pipe_rxsynchd1,              //                   .rxsynchd1
		input  wire [1:0]  hip_pipe_rxsynchd2,              //                   .rxsynchd2
		input  wire [1:0]  hip_pipe_rxsynchd3,              //                   .rxsynchd3
		input  wire [1:0]  hip_pipe_rxsynchd4,              //                   .rxsynchd4
		input  wire [1:0]  hip_pipe_rxsynchd5,              //                   .rxsynchd5
		input  wire [1:0]  hip_pipe_rxsynchd6,              //                   .rxsynchd6
		input  wire [1:0]  hip_pipe_rxsynchd7,              //                   .rxsynchd7
		output wire [17:0] hip_pipe_currentcoeff0,          //                   .currentcoeff0
		output wire [17:0] hip_pipe_currentcoeff1,          //                   .currentcoeff1
		output wire [17:0] hip_pipe_currentcoeff2,          //                   .currentcoeff2
		output wire [17:0] hip_pipe_currentcoeff3,          //                   .currentcoeff3
		output wire [17:0] hip_pipe_currentcoeff4,          //                   .currentcoeff4
		output wire [17:0] hip_pipe_currentcoeff5,          //                   .currentcoeff5
		output wire [17:0] hip_pipe_currentcoeff6,          //                   .currentcoeff6
		output wire [17:0] hip_pipe_currentcoeff7,          //                   .currentcoeff7
		output wire [2:0]  hip_pipe_currentrxpreset0,       //                   .currentrxpreset0
		output wire [2:0]  hip_pipe_currentrxpreset1,       //                   .currentrxpreset1
		output wire [2:0]  hip_pipe_currentrxpreset2,       //                   .currentrxpreset2
		output wire [2:0]  hip_pipe_currentrxpreset3,       //                   .currentrxpreset3
		output wire [2:0]  hip_pipe_currentrxpreset4,       //                   .currentrxpreset4
		output wire [2:0]  hip_pipe_currentrxpreset5,       //                   .currentrxpreset5
		output wire [2:0]  hip_pipe_currentrxpreset6,       //                   .currentrxpreset6
		output wire [2:0]  hip_pipe_currentrxpreset7,       //                   .currentrxpreset7
		output wire [1:0]  hip_pipe_txsynchd0,              //                   .txsynchd0
		output wire [1:0]  hip_pipe_txsynchd1,              //                   .txsynchd1
		output wire [1:0]  hip_pipe_txsynchd2,              //                   .txsynchd2
		output wire [1:0]  hip_pipe_txsynchd3,              //                   .txsynchd3
		output wire [1:0]  hip_pipe_txsynchd4,              //                   .txsynchd4
		output wire [1:0]  hip_pipe_txsynchd5,              //                   .txsynchd5
		output wire [1:0]  hip_pipe_txsynchd6,              //                   .txsynchd6
		output wire [1:0]  hip_pipe_txsynchd7,              //                   .txsynchd7
		output wire        hip_pipe_txblkst0,               //                   .txblkst0
		output wire        hip_pipe_txblkst1,               //                   .txblkst1
		output wire        hip_pipe_txblkst2,               //                   .txblkst2
		output wire        hip_pipe_txblkst3,               //                   .txblkst3
		output wire        hip_pipe_txblkst4,               //                   .txblkst4
		output wire        hip_pipe_txblkst5,               //                   .txblkst5
		output wire        hip_pipe_txblkst6,               //                   .txblkst6
		output wire        hip_pipe_txblkst7,               //                   .txblkst7
		output wire        hip_pipe_txdataskip0,            //                   .txdataskip0
		output wire        hip_pipe_txdataskip1,            //                   .txdataskip1
		output wire        hip_pipe_txdataskip2,            //                   .txdataskip2
		output wire        hip_pipe_txdataskip3,            //                   .txdataskip3
		output wire        hip_pipe_txdataskip4,            //                   .txdataskip4
		output wire        hip_pipe_txdataskip5,            //                   .txdataskip5
		output wire        hip_pipe_txdataskip6,            //                   .txdataskip6
		output wire        hip_pipe_txdataskip7,            //                   .txdataskip7
		output wire [1:0]  hip_pipe_rate0,                  //                   .rate0
		output wire [1:0]  hip_pipe_rate1,                  //                   .rate1
		output wire [1:0]  hip_pipe_rate2,                  //                   .rate2
		output wire [1:0]  hip_pipe_rate3,                  //                   .rate3
		output wire [1:0]  hip_pipe_rate4,                  //                   .rate4
		output wire [1:0]  hip_pipe_rate5,                  //                   .rate5
		output wire [1:0]  hip_pipe_rate6,                  //                   .rate6
		output wire [1:0]  hip_pipe_rate7,                  //                   .rate7
		input  wire        hip_serial_rx_in0,               //         hip_serial.rx_in0
		input  wire        hip_serial_rx_in1,               //                   .rx_in1
		input  wire        hip_serial_rx_in2,               //                   .rx_in2
		input  wire        hip_serial_rx_in3,               //                   .rx_in3
		input  wire        hip_serial_rx_in4,               //                   .rx_in4
		input  wire        hip_serial_rx_in5,               //                   .rx_in5
		input  wire        hip_serial_rx_in6,               //                   .rx_in6
		input  wire        hip_serial_rx_in7,               //                   .rx_in7
		output wire        hip_serial_tx_out0,              //                   .tx_out0
		output wire        hip_serial_tx_out1,              //                   .tx_out1
		output wire        hip_serial_tx_out2,              //                   .tx_out2
		output wire        hip_serial_tx_out3,              //                   .tx_out3
		output wire        hip_serial_tx_out4,              //                   .tx_out4
		output wire        hip_serial_tx_out5,              //                   .tx_out5
		output wire        hip_serial_tx_out6,              //                   .tx_out6
		output wire        hip_serial_tx_out7,              //                   .tx_out7
		input  wire        dut_npor_npor,                   //           dut_npor.npor
		input  wire        dut_npor_pin_perst,              //                   .pin_perst
		input  wire        refclk_clk,                      //             refclk.clk
		output wire        core_clk_out_clk,                //       core_clk_out.clk
		output wire [0:0]  emif_0_mem_mem_ck,               //         emif_0_mem.mem_ck
		output wire [0:0]  emif_0_mem_mem_ck_n,             //                   .mem_ck_n
		output wire [16:0] emif_0_mem_mem_a,                //                   .mem_a
		output wire [0:0]  emif_0_mem_mem_act_n,            //                   .mem_act_n
		output wire [1:0]  emif_0_mem_mem_ba,               //                   .mem_ba
		output wire [0:0]  emif_0_mem_mem_bg,               //                   .mem_bg
		output wire [0:0]  emif_0_mem_mem_cke,              //                   .mem_cke
		output wire [0:0]  emif_0_mem_mem_cs_n,             //                   .mem_cs_n
		output wire [0:0]  emif_0_mem_mem_odt,              //                   .mem_odt
		output wire [0:0]  emif_0_mem_mem_reset_n,          //                   .mem_reset_n
		inout  wire [7:0]  emif_0_mem_mem_dqs,              //                   .mem_dqs
		inout  wire [7:0]  emif_0_mem_mem_dqs_n,            //                   .mem_dqs_n
		inout  wire [63:0] emif_0_mem_mem_dq,               //                   .mem_dq
		inout  wire [7:0]  emif_0_mem_mem_dbi_n,            //                   .mem_dbi_n
		input  wire        emif_0_oct_oct_rzqin,            //         emif_0_oct.oct_rzqin
		input  wire        emif_0_pll_ref_clk_clk,          // emif_0_pll_ref_clk.clk
		output wire        emif_0_status_local_cal_success, //      emif_0_status.local_cal_success
		output wire        emif_0_status_local_cal_fail     //                   .local_cal_fail
	);

	wire          dut_coreclkout_hip_clk;                            // DUT:coreclkout_hip -> [clk_0:in_clk, mm_interconnect_0:DUT_coreclkout_hip_clk, mm_interconnect_1:DUT_coreclkout_hip_clk, onchip_memory2_0:clk, onchip_memory2_0:clk2, rst_controller:clk]
	wire          dut_app_nreset_status_reset;                       // DUT:app_nreset_status -> [clk_0:reset_n, emif_0:global_reset_n, rst_controller:reset_in0]
	wire          dut_dma_rd_master_waitrequest;                     // mm_interconnect_0:DUT_dma_rd_master_waitrequest -> DUT:rd_dma_wait_request_i
	wire   [63:0] dut_dma_rd_master_address;                         // DUT:rd_dma_address_o -> mm_interconnect_0:DUT_dma_rd_master_address
	wire   [31:0] dut_dma_rd_master_byteenable;                      // DUT:rd_dma_byte_enable_o -> mm_interconnect_0:DUT_dma_rd_master_byteenable
	wire          dut_dma_rd_master_write;                           // DUT:rd_dma_write_o -> mm_interconnect_0:DUT_dma_rd_master_write
	wire  [255:0] dut_dma_rd_master_writedata;                       // DUT:rd_dma_write_data_o -> mm_interconnect_0:DUT_dma_rd_master_writedata
	wire    [4:0] dut_dma_rd_master_burstcount;                      // DUT:rd_dma_burst_count_o -> mm_interconnect_0:DUT_dma_rd_master_burstcount
	wire  [255:0] dut_dma_wr_master_readdata;                        // mm_interconnect_0:DUT_dma_wr_master_readdata -> DUT:wr_dma_read_data_i
	wire          dut_dma_wr_master_waitrequest;                     // mm_interconnect_0:DUT_dma_wr_master_waitrequest -> DUT:wr_dma_wait_request_i
	wire   [63:0] dut_dma_wr_master_address;                         // DUT:wr_dma_address_o -> mm_interconnect_0:DUT_dma_wr_master_address
	wire          dut_dma_wr_master_read;                            // DUT:wr_dma_read_o -> mm_interconnect_0:DUT_dma_wr_master_read
	wire          dut_dma_wr_master_readdatavalid;                   // mm_interconnect_0:DUT_dma_wr_master_readdatavalid -> DUT:wr_dma_read_data_valid_i
	wire    [4:0] dut_dma_wr_master_burstcount;                      // DUT:wr_dma_burst_count_o -> mm_interconnect_0:DUT_dma_wr_master_burstcount
	wire   [31:0] dut_rxm_bar2_readdata;                             // mm_interconnect_0:DUT_rxm_bar2_readdata -> DUT:rxm_bar2_readdata_i
	wire          dut_rxm_bar2_waitrequest;                          // mm_interconnect_0:DUT_rxm_bar2_waitrequest -> DUT:rxm_bar2_waitrequest_i
	wire   [63:0] dut_rxm_bar2_address;                              // DUT:rxm_bar2_address_o -> mm_interconnect_0:DUT_rxm_bar2_address
	wire    [3:0] dut_rxm_bar2_byteenable;                           // DUT:rxm_bar2_byteenable_o -> mm_interconnect_0:DUT_rxm_bar2_byteenable
	wire          dut_rxm_bar2_read;                                 // DUT:rxm_bar2_read_o -> mm_interconnect_0:DUT_rxm_bar2_read
	wire          dut_rxm_bar2_readdatavalid;                        // mm_interconnect_0:DUT_rxm_bar2_readdatavalid -> DUT:rxm_bar2_readdatavalid_i
	wire   [31:0] dut_rxm_bar2_writedata;                            // DUT:rxm_bar2_writedata_o -> mm_interconnect_0:DUT_rxm_bar2_writedata
	wire          dut_rxm_bar2_write;                                // DUT:rxm_bar2_write_o -> mm_interconnect_0:DUT_rxm_bar2_write
	wire  [511:0] mm_interconnect_0_emif_0_ctrl_amm_0_readdata;      // emif_0:amm_readdata_0 -> mm_interconnect_0:emif_0_ctrl_amm_0_readdata
	wire          mm_interconnect_0_emif_0_ctrl_amm_0_waitrequest;   // emif_0:amm_ready_0 -> mm_interconnect_0:emif_0_ctrl_amm_0_waitrequest
	wire   [21:0] mm_interconnect_0_emif_0_ctrl_amm_0_address;       // mm_interconnect_0:emif_0_ctrl_amm_0_address -> emif_0:amm_address_0
	wire          mm_interconnect_0_emif_0_ctrl_amm_0_read;          // mm_interconnect_0:emif_0_ctrl_amm_0_read -> emif_0:amm_read_0
	wire   [63:0] mm_interconnect_0_emif_0_ctrl_amm_0_byteenable;    // mm_interconnect_0:emif_0_ctrl_amm_0_byteenable -> emif_0:amm_byteenable_0
	wire          mm_interconnect_0_emif_0_ctrl_amm_0_readdatavalid; // emif_0:amm_readdatavalid_0 -> mm_interconnect_0:emif_0_ctrl_amm_0_readdatavalid
	wire          mm_interconnect_0_emif_0_ctrl_amm_0_write;         // mm_interconnect_0:emif_0_ctrl_amm_0_write -> emif_0:amm_write_0
	wire  [511:0] mm_interconnect_0_emif_0_ctrl_amm_0_writedata;     // mm_interconnect_0:emif_0_ctrl_amm_0_writedata -> emif_0:amm_writedata_0
	wire    [6:0] mm_interconnect_0_emif_0_ctrl_amm_0_burstcount;    // mm_interconnect_0:emif_0_ctrl_amm_0_burstcount -> emif_0:amm_burstcount_0
	wire          emif_0_emif_usr_clk_clk;                           // emif_0:emif_usr_clk -> [mm_interconnect_0:emif_0_emif_usr_clk_clk, rst_controller_001:clk]
	wire          mm_interconnect_0_dut_rd_dts_slave_chipselect;     // mm_interconnect_0:DUT_rd_dts_slave_chipselect -> DUT:rd_dts_chip_select_i
	wire          mm_interconnect_0_dut_rd_dts_slave_waitrequest;    // DUT:rd_dts_wait_request_o -> mm_interconnect_0:DUT_rd_dts_slave_waitrequest
	wire    [7:0] mm_interconnect_0_dut_rd_dts_slave_address;        // mm_interconnect_0:DUT_rd_dts_slave_address -> DUT:rd_dts_address_i
	wire          mm_interconnect_0_dut_rd_dts_slave_write;          // mm_interconnect_0:DUT_rd_dts_slave_write -> DUT:rd_dts_write_i
	wire  [255:0] mm_interconnect_0_dut_rd_dts_slave_writedata;      // mm_interconnect_0:DUT_rd_dts_slave_writedata -> DUT:rd_dts_write_data_i
	wire    [4:0] mm_interconnect_0_dut_rd_dts_slave_burstcount;     // mm_interconnect_0:DUT_rd_dts_slave_burstcount -> DUT:rd_dts_burst_count_i
	wire          mm_interconnect_0_onchip_memory2_0_s2_chipselect;  // mm_interconnect_0:onchip_memory2_0_s2_chipselect -> onchip_memory2_0:chipselect2
	wire  [255:0] mm_interconnect_0_onchip_memory2_0_s2_readdata;    // onchip_memory2_0:readdata2 -> mm_interconnect_0:onchip_memory2_0_s2_readdata
	wire   [10:0] mm_interconnect_0_onchip_memory2_0_s2_address;     // mm_interconnect_0:onchip_memory2_0_s2_address -> onchip_memory2_0:address2
	wire   [31:0] mm_interconnect_0_onchip_memory2_0_s2_byteenable;  // mm_interconnect_0:onchip_memory2_0_s2_byteenable -> onchip_memory2_0:byteenable2
	wire          mm_interconnect_0_onchip_memory2_0_s2_write;       // mm_interconnect_0:onchip_memory2_0_s2_write -> onchip_memory2_0:write2
	wire  [255:0] mm_interconnect_0_onchip_memory2_0_s2_writedata;   // mm_interconnect_0:onchip_memory2_0_s2_writedata -> onchip_memory2_0:writedata2
	wire          mm_interconnect_0_onchip_memory2_0_s2_clken;       // mm_interconnect_0:onchip_memory2_0_s2_clken -> onchip_memory2_0:clken2
	wire          mm_interconnect_0_dut_wr_dts_slave_chipselect;     // mm_interconnect_0:DUT_wr_dts_slave_chipselect -> DUT:wr_dts_chip_select_i
	wire          mm_interconnect_0_dut_wr_dts_slave_waitrequest;    // DUT:wr_dts_wait_request_o -> mm_interconnect_0:DUT_wr_dts_slave_waitrequest
	wire    [7:0] mm_interconnect_0_dut_wr_dts_slave_address;        // mm_interconnect_0:DUT_wr_dts_slave_address -> DUT:wr_dts_address_i
	wire          mm_interconnect_0_dut_wr_dts_slave_write;          // mm_interconnect_0:DUT_wr_dts_slave_write -> DUT:wr_dts_write_i
	wire  [255:0] mm_interconnect_0_dut_wr_dts_slave_writedata;      // mm_interconnect_0:DUT_wr_dts_slave_writedata -> DUT:wr_dts_write_data_i
	wire    [4:0] mm_interconnect_0_dut_wr_dts_slave_burstcount;     // mm_interconnect_0:DUT_wr_dts_slave_burstcount -> DUT:wr_dts_burst_count_i
	wire          mm_interconnect_0_onchip_memory2_0_s1_chipselect;  // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [255:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;    // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [10:0] mm_interconnect_0_onchip_memory2_0_s1_address;     // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [31:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;  // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire          mm_interconnect_0_onchip_memory2_0_s1_write;       // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [255:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;   // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire          mm_interconnect_0_onchip_memory2_0_s1_clken;       // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire          dut_rd_dcm_master_waitrequest;                     // mm_interconnect_1:DUT_rd_dcm_master_waitrequest -> DUT:rd_dcm_wait_request_i
	wire   [31:0] dut_rd_dcm_master_readdata;                        // mm_interconnect_1:DUT_rd_dcm_master_readdata -> DUT:rd_dcm_read_data_i
	wire   [63:0] dut_rd_dcm_master_address;                         // DUT:rd_dcm_address_o -> mm_interconnect_1:DUT_rd_dcm_master_address
	wire          dut_rd_dcm_master_read;                            // DUT:rd_dcm_read_o -> mm_interconnect_1:DUT_rd_dcm_master_read
	wire    [3:0] dut_rd_dcm_master_byteenable;                      // DUT:rd_dcm_byte_enable_o -> mm_interconnect_1:DUT_rd_dcm_master_byteenable
	wire          dut_rd_dcm_master_readdatavalid;                   // mm_interconnect_1:DUT_rd_dcm_master_readdatavalid -> DUT:rd_dcm_read_data_valid_i
	wire          dut_rd_dcm_master_write;                           // DUT:rd_dcm_write_o -> mm_interconnect_1:DUT_rd_dcm_master_write
	wire   [31:0] dut_rd_dcm_master_writedata;                       // DUT:rd_dcm_writedata_o -> mm_interconnect_1:DUT_rd_dcm_master_writedata
	wire          dut_wr_dcm_master_waitrequest;                     // mm_interconnect_1:DUT_wr_dcm_master_waitrequest -> DUT:wr_dcm_wait_request_i
	wire   [31:0] dut_wr_dcm_master_readdata;                        // mm_interconnect_1:DUT_wr_dcm_master_readdata -> DUT:wr_dcm_read_data_i
	wire   [63:0] dut_wr_dcm_master_address;                         // DUT:wr_dcm_address_o -> mm_interconnect_1:DUT_wr_dcm_master_address
	wire          dut_wr_dcm_master_read;                            // DUT:wr_dcm_read_o -> mm_interconnect_1:DUT_wr_dcm_master_read
	wire    [3:0] dut_wr_dcm_master_byteenable;                      // DUT:wr_dcm_byte_enable_o -> mm_interconnect_1:DUT_wr_dcm_master_byteenable
	wire          dut_wr_dcm_master_readdatavalid;                   // mm_interconnect_1:DUT_wr_dcm_master_readdatavalid -> DUT:wr_dcm_read_data_valid_i
	wire          dut_wr_dcm_master_write;                           // DUT:wr_dcm_write_o -> mm_interconnect_1:DUT_wr_dcm_master_write
	wire   [31:0] dut_wr_dcm_master_writedata;                       // DUT:wr_dcm_writedata_o -> mm_interconnect_1:DUT_wr_dcm_master_writedata
	wire          mm_interconnect_1_dut_txs_chipselect;              // mm_interconnect_1:DUT_txs_chipselect -> DUT:txs_chipselect_i
	wire   [31:0] mm_interconnect_1_dut_txs_readdata;                // DUT:txs_readdata_o -> mm_interconnect_1:DUT_txs_readdata
	wire          mm_interconnect_1_dut_txs_waitrequest;             // DUT:txs_waitrequest_o -> mm_interconnect_1:DUT_txs_waitrequest
	wire   [39:0] mm_interconnect_1_dut_txs_address;                 // mm_interconnect_1:DUT_txs_address -> DUT:txs_address_i
	wire          mm_interconnect_1_dut_txs_read;                    // mm_interconnect_1:DUT_txs_read -> DUT:txs_read_i
	wire    [3:0] mm_interconnect_1_dut_txs_byteenable;              // mm_interconnect_1:DUT_txs_byteenable -> DUT:txs_byteenable_i
	wire          mm_interconnect_1_dut_txs_readdatavalid;           // DUT:txs_readdatavalid_o -> mm_interconnect_1:DUT_txs_readdatavalid
	wire          mm_interconnect_1_dut_txs_write;                   // mm_interconnect_1:DUT_txs_write -> DUT:txs_write_i
	wire   [31:0] mm_interconnect_1_dut_txs_writedata;               // mm_interconnect_1:DUT_txs_writedata -> DUT:txs_writedata_i
	wire          rst_controller_reset_out_reset;                    // rst_controller:reset_out -> [mm_interconnect_0:onchip_memory2_0_reset2_reset_bridge_in_reset_reset, mm_interconnect_1:DUT_rd_dcm_master_translator_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, onchip_memory2_0:reset2]
	wire          rst_controller_reset_out_reset_req;                // rst_controller:reset_req -> [onchip_memory2_0:reset_req, onchip_memory2_0:reset_req2, rst_translator:reset_req_in]
	wire          rst_controller_001_reset_out_reset;                // rst_controller_001:reset_out -> mm_interconnect_0:emif_0_ctrl_amm_0_translator_reset_reset_bridge_in_reset_reset
	wire          emif_0_emif_usr_reset_n_reset;                     // emif_0:emif_usr_reset_n -> rst_controller_001:reset_in0

	top_DUT dut (
		.app_nreset_status        (dut_app_nreset_status_reset),                    //  output,    width = 1, app_nreset_status.reset_n
		.coreclkout_hip           (dut_coreclkout_hip_clk),                         //  output,    width = 1,    coreclkout_hip.clk
		.rd_dma_address_o         (dut_dma_rd_master_address),                      //  output,   width = 64,     dma_rd_master.address
		.rd_dma_write_o           (dut_dma_rd_master_write),                        //  output,    width = 1,                  .write
		.rd_dma_write_data_o      (dut_dma_rd_master_writedata),                    //  output,  width = 256,                  .writedata
		.rd_dma_wait_request_i    (dut_dma_rd_master_waitrequest),                  //   input,    width = 1,                  .waitrequest
		.rd_dma_burst_count_o     (dut_dma_rd_master_burstcount),                   //  output,    width = 5,                  .burstcount
		.rd_dma_byte_enable_o     (dut_dma_rd_master_byteenable),                   //  output,   width = 32,                  .byteenable
		.wr_dma_address_o         (dut_dma_wr_master_address),                      //  output,   width = 64,     dma_wr_master.address
		.wr_dma_read_o            (dut_dma_wr_master_read),                         //  output,    width = 1,                  .read
		.wr_dma_read_data_i       (dut_dma_wr_master_readdata),                     //   input,  width = 256,                  .readdata
		.wr_dma_wait_request_i    (dut_dma_wr_master_waitrequest),                  //   input,    width = 1,                  .waitrequest
		.wr_dma_burst_count_o     (dut_dma_wr_master_burstcount),                   //  output,    width = 5,                  .burstcount
		.wr_dma_read_data_valid_i (dut_dma_wr_master_readdatavalid),                //   input,    width = 1,                  .readdatavalid
		.test_in                  (hip_ctrl_test_in),                               //   input,   width = 32,          hip_ctrl.test_in
		.simu_mode_pipe           (hip_ctrl_simu_mode_pipe),                        //   input,    width = 1,                  .simu_mode_pipe
		.sim_pipe_pclk_in         (hip_pipe_sim_pipe_pclk_in),                      //   input,    width = 1,          hip_pipe.sim_pipe_pclk_in
		.sim_pipe_rate            (hip_pipe_sim_pipe_rate),                         //  output,    width = 2,                  .sim_pipe_rate
		.sim_ltssmstate           (hip_pipe_sim_ltssmstate),                        //  output,    width = 5,                  .sim_ltssmstate
		.eidleinfersel0           (hip_pipe_eidleinfersel0),                        //  output,    width = 3,                  .eidleinfersel0
		.eidleinfersel1           (hip_pipe_eidleinfersel1),                        //  output,    width = 3,                  .eidleinfersel1
		.eidleinfersel2           (hip_pipe_eidleinfersel2),                        //  output,    width = 3,                  .eidleinfersel2
		.eidleinfersel3           (hip_pipe_eidleinfersel3),                        //  output,    width = 3,                  .eidleinfersel3
		.eidleinfersel4           (hip_pipe_eidleinfersel4),                        //  output,    width = 3,                  .eidleinfersel4
		.eidleinfersel5           (hip_pipe_eidleinfersel5),                        //  output,    width = 3,                  .eidleinfersel5
		.eidleinfersel6           (hip_pipe_eidleinfersel6),                        //  output,    width = 3,                  .eidleinfersel6
		.eidleinfersel7           (hip_pipe_eidleinfersel7),                        //  output,    width = 3,                  .eidleinfersel7
		.powerdown0               (hip_pipe_powerdown0),                            //  output,    width = 2,                  .powerdown0
		.powerdown1               (hip_pipe_powerdown1),                            //  output,    width = 2,                  .powerdown1
		.powerdown2               (hip_pipe_powerdown2),                            //  output,    width = 2,                  .powerdown2
		.powerdown3               (hip_pipe_powerdown3),                            //  output,    width = 2,                  .powerdown3
		.powerdown4               (hip_pipe_powerdown4),                            //  output,    width = 2,                  .powerdown4
		.powerdown5               (hip_pipe_powerdown5),                            //  output,    width = 2,                  .powerdown5
		.powerdown6               (hip_pipe_powerdown6),                            //  output,    width = 2,                  .powerdown6
		.powerdown7               (hip_pipe_powerdown7),                            //  output,    width = 2,                  .powerdown7
		.rxpolarity0              (hip_pipe_rxpolarity0),                           //  output,    width = 1,                  .rxpolarity0
		.rxpolarity1              (hip_pipe_rxpolarity1),                           //  output,    width = 1,                  .rxpolarity1
		.rxpolarity2              (hip_pipe_rxpolarity2),                           //  output,    width = 1,                  .rxpolarity2
		.rxpolarity3              (hip_pipe_rxpolarity3),                           //  output,    width = 1,                  .rxpolarity3
		.rxpolarity4              (hip_pipe_rxpolarity4),                           //  output,    width = 1,                  .rxpolarity4
		.rxpolarity5              (hip_pipe_rxpolarity5),                           //  output,    width = 1,                  .rxpolarity5
		.rxpolarity6              (hip_pipe_rxpolarity6),                           //  output,    width = 1,                  .rxpolarity6
		.rxpolarity7              (hip_pipe_rxpolarity7),                           //  output,    width = 1,                  .rxpolarity7
		.txcompl0                 (hip_pipe_txcompl0),                              //  output,    width = 1,                  .txcompl0
		.txcompl1                 (hip_pipe_txcompl1),                              //  output,    width = 1,                  .txcompl1
		.txcompl2                 (hip_pipe_txcompl2),                              //  output,    width = 1,                  .txcompl2
		.txcompl3                 (hip_pipe_txcompl3),                              //  output,    width = 1,                  .txcompl3
		.txcompl4                 (hip_pipe_txcompl4),                              //  output,    width = 1,                  .txcompl4
		.txcompl5                 (hip_pipe_txcompl5),                              //  output,    width = 1,                  .txcompl5
		.txcompl6                 (hip_pipe_txcompl6),                              //  output,    width = 1,                  .txcompl6
		.txcompl7                 (hip_pipe_txcompl7),                              //  output,    width = 1,                  .txcompl7
		.txdata0                  (hip_pipe_txdata0),                               //  output,   width = 32,                  .txdata0
		.txdata1                  (hip_pipe_txdata1),                               //  output,   width = 32,                  .txdata1
		.txdata2                  (hip_pipe_txdata2),                               //  output,   width = 32,                  .txdata2
		.txdata3                  (hip_pipe_txdata3),                               //  output,   width = 32,                  .txdata3
		.txdata4                  (hip_pipe_txdata4),                               //  output,   width = 32,                  .txdata4
		.txdata5                  (hip_pipe_txdata5),                               //  output,   width = 32,                  .txdata5
		.txdata6                  (hip_pipe_txdata6),                               //  output,   width = 32,                  .txdata6
		.txdata7                  (hip_pipe_txdata7),                               //  output,   width = 32,                  .txdata7
		.txdatak0                 (hip_pipe_txdatak0),                              //  output,    width = 4,                  .txdatak0
		.txdatak1                 (hip_pipe_txdatak1),                              //  output,    width = 4,                  .txdatak1
		.txdatak2                 (hip_pipe_txdatak2),                              //  output,    width = 4,                  .txdatak2
		.txdatak3                 (hip_pipe_txdatak3),                              //  output,    width = 4,                  .txdatak3
		.txdatak4                 (hip_pipe_txdatak4),                              //  output,    width = 4,                  .txdatak4
		.txdatak5                 (hip_pipe_txdatak5),                              //  output,    width = 4,                  .txdatak5
		.txdatak6                 (hip_pipe_txdatak6),                              //  output,    width = 4,                  .txdatak6
		.txdatak7                 (hip_pipe_txdatak7),                              //  output,    width = 4,                  .txdatak7
		.txdetectrx0              (hip_pipe_txdetectrx0),                           //  output,    width = 1,                  .txdetectrx0
		.txdetectrx1              (hip_pipe_txdetectrx1),                           //  output,    width = 1,                  .txdetectrx1
		.txdetectrx2              (hip_pipe_txdetectrx2),                           //  output,    width = 1,                  .txdetectrx2
		.txdetectrx3              (hip_pipe_txdetectrx3),                           //  output,    width = 1,                  .txdetectrx3
		.txdetectrx4              (hip_pipe_txdetectrx4),                           //  output,    width = 1,                  .txdetectrx4
		.txdetectrx5              (hip_pipe_txdetectrx5),                           //  output,    width = 1,                  .txdetectrx5
		.txdetectrx6              (hip_pipe_txdetectrx6),                           //  output,    width = 1,                  .txdetectrx6
		.txdetectrx7              (hip_pipe_txdetectrx7),                           //  output,    width = 1,                  .txdetectrx7
		.txelecidle0              (hip_pipe_txelecidle0),                           //  output,    width = 1,                  .txelecidle0
		.txelecidle1              (hip_pipe_txelecidle1),                           //  output,    width = 1,                  .txelecidle1
		.txelecidle2              (hip_pipe_txelecidle2),                           //  output,    width = 1,                  .txelecidle2
		.txelecidle3              (hip_pipe_txelecidle3),                           //  output,    width = 1,                  .txelecidle3
		.txelecidle4              (hip_pipe_txelecidle4),                           //  output,    width = 1,                  .txelecidle4
		.txelecidle5              (hip_pipe_txelecidle5),                           //  output,    width = 1,                  .txelecidle5
		.txelecidle6              (hip_pipe_txelecidle6),                           //  output,    width = 1,                  .txelecidle6
		.txelecidle7              (hip_pipe_txelecidle7),                           //  output,    width = 1,                  .txelecidle7
		.txdeemph0                (hip_pipe_txdeemph0),                             //  output,    width = 1,                  .txdeemph0
		.txdeemph1                (hip_pipe_txdeemph1),                             //  output,    width = 1,                  .txdeemph1
		.txdeemph2                (hip_pipe_txdeemph2),                             //  output,    width = 1,                  .txdeemph2
		.txdeemph3                (hip_pipe_txdeemph3),                             //  output,    width = 1,                  .txdeemph3
		.txdeemph4                (hip_pipe_txdeemph4),                             //  output,    width = 1,                  .txdeemph4
		.txdeemph5                (hip_pipe_txdeemph5),                             //  output,    width = 1,                  .txdeemph5
		.txdeemph6                (hip_pipe_txdeemph6),                             //  output,    width = 1,                  .txdeemph6
		.txdeemph7                (hip_pipe_txdeemph7),                             //  output,    width = 1,                  .txdeemph7
		.txmargin0                (hip_pipe_txmargin0),                             //  output,    width = 3,                  .txmargin0
		.txmargin1                (hip_pipe_txmargin1),                             //  output,    width = 3,                  .txmargin1
		.txmargin2                (hip_pipe_txmargin2),                             //  output,    width = 3,                  .txmargin2
		.txmargin3                (hip_pipe_txmargin3),                             //  output,    width = 3,                  .txmargin3
		.txmargin4                (hip_pipe_txmargin4),                             //  output,    width = 3,                  .txmargin4
		.txmargin5                (hip_pipe_txmargin5),                             //  output,    width = 3,                  .txmargin5
		.txmargin6                (hip_pipe_txmargin6),                             //  output,    width = 3,                  .txmargin6
		.txmargin7                (hip_pipe_txmargin7),                             //  output,    width = 3,                  .txmargin7
		.txswing0                 (hip_pipe_txswing0),                              //  output,    width = 1,                  .txswing0
		.txswing1                 (hip_pipe_txswing1),                              //  output,    width = 1,                  .txswing1
		.txswing2                 (hip_pipe_txswing2),                              //  output,    width = 1,                  .txswing2
		.txswing3                 (hip_pipe_txswing3),                              //  output,    width = 1,                  .txswing3
		.txswing4                 (hip_pipe_txswing4),                              //  output,    width = 1,                  .txswing4
		.txswing5                 (hip_pipe_txswing5),                              //  output,    width = 1,                  .txswing5
		.txswing6                 (hip_pipe_txswing6),                              //  output,    width = 1,                  .txswing6
		.txswing7                 (hip_pipe_txswing7),                              //  output,    width = 1,                  .txswing7
		.phystatus0               (hip_pipe_phystatus0),                            //   input,    width = 1,                  .phystatus0
		.phystatus1               (hip_pipe_phystatus1),                            //   input,    width = 1,                  .phystatus1
		.phystatus2               (hip_pipe_phystatus2),                            //   input,    width = 1,                  .phystatus2
		.phystatus3               (hip_pipe_phystatus3),                            //   input,    width = 1,                  .phystatus3
		.phystatus4               (hip_pipe_phystatus4),                            //   input,    width = 1,                  .phystatus4
		.phystatus5               (hip_pipe_phystatus5),                            //   input,    width = 1,                  .phystatus5
		.phystatus6               (hip_pipe_phystatus6),                            //   input,    width = 1,                  .phystatus6
		.phystatus7               (hip_pipe_phystatus7),                            //   input,    width = 1,                  .phystatus7
		.rxdata0                  (hip_pipe_rxdata0),                               //   input,   width = 32,                  .rxdata0
		.rxdata1                  (hip_pipe_rxdata1),                               //   input,   width = 32,                  .rxdata1
		.rxdata2                  (hip_pipe_rxdata2),                               //   input,   width = 32,                  .rxdata2
		.rxdata3                  (hip_pipe_rxdata3),                               //   input,   width = 32,                  .rxdata3
		.rxdata4                  (hip_pipe_rxdata4),                               //   input,   width = 32,                  .rxdata4
		.rxdata5                  (hip_pipe_rxdata5),                               //   input,   width = 32,                  .rxdata5
		.rxdata6                  (hip_pipe_rxdata6),                               //   input,   width = 32,                  .rxdata6
		.rxdata7                  (hip_pipe_rxdata7),                               //   input,   width = 32,                  .rxdata7
		.rxdatak0                 (hip_pipe_rxdatak0),                              //   input,    width = 4,                  .rxdatak0
		.rxdatak1                 (hip_pipe_rxdatak1),                              //   input,    width = 4,                  .rxdatak1
		.rxdatak2                 (hip_pipe_rxdatak2),                              //   input,    width = 4,                  .rxdatak2
		.rxdatak3                 (hip_pipe_rxdatak3),                              //   input,    width = 4,                  .rxdatak3
		.rxdatak4                 (hip_pipe_rxdatak4),                              //   input,    width = 4,                  .rxdatak4
		.rxdatak5                 (hip_pipe_rxdatak5),                              //   input,    width = 4,                  .rxdatak5
		.rxdatak6                 (hip_pipe_rxdatak6),                              //   input,    width = 4,                  .rxdatak6
		.rxdatak7                 (hip_pipe_rxdatak7),                              //   input,    width = 4,                  .rxdatak7
		.rxelecidle0              (hip_pipe_rxelecidle0),                           //   input,    width = 1,                  .rxelecidle0
		.rxelecidle1              (hip_pipe_rxelecidle1),                           //   input,    width = 1,                  .rxelecidle1
		.rxelecidle2              (hip_pipe_rxelecidle2),                           //   input,    width = 1,                  .rxelecidle2
		.rxelecidle3              (hip_pipe_rxelecidle3),                           //   input,    width = 1,                  .rxelecidle3
		.rxelecidle4              (hip_pipe_rxelecidle4),                           //   input,    width = 1,                  .rxelecidle4
		.rxelecidle5              (hip_pipe_rxelecidle5),                           //   input,    width = 1,                  .rxelecidle5
		.rxelecidle6              (hip_pipe_rxelecidle6),                           //   input,    width = 1,                  .rxelecidle6
		.rxelecidle7              (hip_pipe_rxelecidle7),                           //   input,    width = 1,                  .rxelecidle7
		.rxstatus0                (hip_pipe_rxstatus0),                             //   input,    width = 3,                  .rxstatus0
		.rxstatus1                (hip_pipe_rxstatus1),                             //   input,    width = 3,                  .rxstatus1
		.rxstatus2                (hip_pipe_rxstatus2),                             //   input,    width = 3,                  .rxstatus2
		.rxstatus3                (hip_pipe_rxstatus3),                             //   input,    width = 3,                  .rxstatus3
		.rxstatus4                (hip_pipe_rxstatus4),                             //   input,    width = 3,                  .rxstatus4
		.rxstatus5                (hip_pipe_rxstatus5),                             //   input,    width = 3,                  .rxstatus5
		.rxstatus6                (hip_pipe_rxstatus6),                             //   input,    width = 3,                  .rxstatus6
		.rxstatus7                (hip_pipe_rxstatus7),                             //   input,    width = 3,                  .rxstatus7
		.rxvalid0                 (hip_pipe_rxvalid0),                              //   input,    width = 1,                  .rxvalid0
		.rxvalid1                 (hip_pipe_rxvalid1),                              //   input,    width = 1,                  .rxvalid1
		.rxvalid2                 (hip_pipe_rxvalid2),                              //   input,    width = 1,                  .rxvalid2
		.rxvalid3                 (hip_pipe_rxvalid3),                              //   input,    width = 1,                  .rxvalid3
		.rxvalid4                 (hip_pipe_rxvalid4),                              //   input,    width = 1,                  .rxvalid4
		.rxvalid5                 (hip_pipe_rxvalid5),                              //   input,    width = 1,                  .rxvalid5
		.rxvalid6                 (hip_pipe_rxvalid6),                              //   input,    width = 1,                  .rxvalid6
		.rxvalid7                 (hip_pipe_rxvalid7),                              //   input,    width = 1,                  .rxvalid7
		.rxdataskip0              (hip_pipe_rxdataskip0),                           //   input,    width = 1,                  .rxdataskip0
		.rxdataskip1              (hip_pipe_rxdataskip1),                           //   input,    width = 1,                  .rxdataskip1
		.rxdataskip2              (hip_pipe_rxdataskip2),                           //   input,    width = 1,                  .rxdataskip2
		.rxdataskip3              (hip_pipe_rxdataskip3),                           //   input,    width = 1,                  .rxdataskip3
		.rxdataskip4              (hip_pipe_rxdataskip4),                           //   input,    width = 1,                  .rxdataskip4
		.rxdataskip5              (hip_pipe_rxdataskip5),                           //   input,    width = 1,                  .rxdataskip5
		.rxdataskip6              (hip_pipe_rxdataskip6),                           //   input,    width = 1,                  .rxdataskip6
		.rxdataskip7              (hip_pipe_rxdataskip7),                           //   input,    width = 1,                  .rxdataskip7
		.rxblkst0                 (hip_pipe_rxblkst0),                              //   input,    width = 1,                  .rxblkst0
		.rxblkst1                 (hip_pipe_rxblkst1),                              //   input,    width = 1,                  .rxblkst1
		.rxblkst2                 (hip_pipe_rxblkst2),                              //   input,    width = 1,                  .rxblkst2
		.rxblkst3                 (hip_pipe_rxblkst3),                              //   input,    width = 1,                  .rxblkst3
		.rxblkst4                 (hip_pipe_rxblkst4),                              //   input,    width = 1,                  .rxblkst4
		.rxblkst5                 (hip_pipe_rxblkst5),                              //   input,    width = 1,                  .rxblkst5
		.rxblkst6                 (hip_pipe_rxblkst6),                              //   input,    width = 1,                  .rxblkst6
		.rxblkst7                 (hip_pipe_rxblkst7),                              //   input,    width = 1,                  .rxblkst7
		.rxsynchd0                (hip_pipe_rxsynchd0),                             //   input,    width = 2,                  .rxsynchd0
		.rxsynchd1                (hip_pipe_rxsynchd1),                             //   input,    width = 2,                  .rxsynchd1
		.rxsynchd2                (hip_pipe_rxsynchd2),                             //   input,    width = 2,                  .rxsynchd2
		.rxsynchd3                (hip_pipe_rxsynchd3),                             //   input,    width = 2,                  .rxsynchd3
		.rxsynchd4                (hip_pipe_rxsynchd4),                             //   input,    width = 2,                  .rxsynchd4
		.rxsynchd5                (hip_pipe_rxsynchd5),                             //   input,    width = 2,                  .rxsynchd5
		.rxsynchd6                (hip_pipe_rxsynchd6),                             //   input,    width = 2,                  .rxsynchd6
		.rxsynchd7                (hip_pipe_rxsynchd7),                             //   input,    width = 2,                  .rxsynchd7
		.currentcoeff0            (hip_pipe_currentcoeff0),                         //  output,   width = 18,                  .currentcoeff0
		.currentcoeff1            (hip_pipe_currentcoeff1),                         //  output,   width = 18,                  .currentcoeff1
		.currentcoeff2            (hip_pipe_currentcoeff2),                         //  output,   width = 18,                  .currentcoeff2
		.currentcoeff3            (hip_pipe_currentcoeff3),                         //  output,   width = 18,                  .currentcoeff3
		.currentcoeff4            (hip_pipe_currentcoeff4),                         //  output,   width = 18,                  .currentcoeff4
		.currentcoeff5            (hip_pipe_currentcoeff5),                         //  output,   width = 18,                  .currentcoeff5
		.currentcoeff6            (hip_pipe_currentcoeff6),                         //  output,   width = 18,                  .currentcoeff6
		.currentcoeff7            (hip_pipe_currentcoeff7),                         //  output,   width = 18,                  .currentcoeff7
		.currentrxpreset0         (hip_pipe_currentrxpreset0),                      //  output,    width = 3,                  .currentrxpreset0
		.currentrxpreset1         (hip_pipe_currentrxpreset1),                      //  output,    width = 3,                  .currentrxpreset1
		.currentrxpreset2         (hip_pipe_currentrxpreset2),                      //  output,    width = 3,                  .currentrxpreset2
		.currentrxpreset3         (hip_pipe_currentrxpreset3),                      //  output,    width = 3,                  .currentrxpreset3
		.currentrxpreset4         (hip_pipe_currentrxpreset4),                      //  output,    width = 3,                  .currentrxpreset4
		.currentrxpreset5         (hip_pipe_currentrxpreset5),                      //  output,    width = 3,                  .currentrxpreset5
		.currentrxpreset6         (hip_pipe_currentrxpreset6),                      //  output,    width = 3,                  .currentrxpreset6
		.currentrxpreset7         (hip_pipe_currentrxpreset7),                      //  output,    width = 3,                  .currentrxpreset7
		.txsynchd0                (hip_pipe_txsynchd0),                             //  output,    width = 2,                  .txsynchd0
		.txsynchd1                (hip_pipe_txsynchd1),                             //  output,    width = 2,                  .txsynchd1
		.txsynchd2                (hip_pipe_txsynchd2),                             //  output,    width = 2,                  .txsynchd2
		.txsynchd3                (hip_pipe_txsynchd3),                             //  output,    width = 2,                  .txsynchd3
		.txsynchd4                (hip_pipe_txsynchd4),                             //  output,    width = 2,                  .txsynchd4
		.txsynchd5                (hip_pipe_txsynchd5),                             //  output,    width = 2,                  .txsynchd5
		.txsynchd6                (hip_pipe_txsynchd6),                             //  output,    width = 2,                  .txsynchd6
		.txsynchd7                (hip_pipe_txsynchd7),                             //  output,    width = 2,                  .txsynchd7
		.txblkst0                 (hip_pipe_txblkst0),                              //  output,    width = 1,                  .txblkst0
		.txblkst1                 (hip_pipe_txblkst1),                              //  output,    width = 1,                  .txblkst1
		.txblkst2                 (hip_pipe_txblkst2),                              //  output,    width = 1,                  .txblkst2
		.txblkst3                 (hip_pipe_txblkst3),                              //  output,    width = 1,                  .txblkst3
		.txblkst4                 (hip_pipe_txblkst4),                              //  output,    width = 1,                  .txblkst4
		.txblkst5                 (hip_pipe_txblkst5),                              //  output,    width = 1,                  .txblkst5
		.txblkst6                 (hip_pipe_txblkst6),                              //  output,    width = 1,                  .txblkst6
		.txblkst7                 (hip_pipe_txblkst7),                              //  output,    width = 1,                  .txblkst7
		.txdataskip0              (hip_pipe_txdataskip0),                           //  output,    width = 1,                  .txdataskip0
		.txdataskip1              (hip_pipe_txdataskip1),                           //  output,    width = 1,                  .txdataskip1
		.txdataskip2              (hip_pipe_txdataskip2),                           //  output,    width = 1,                  .txdataskip2
		.txdataskip3              (hip_pipe_txdataskip3),                           //  output,    width = 1,                  .txdataskip3
		.txdataskip4              (hip_pipe_txdataskip4),                           //  output,    width = 1,                  .txdataskip4
		.txdataskip5              (hip_pipe_txdataskip5),                           //  output,    width = 1,                  .txdataskip5
		.txdataskip6              (hip_pipe_txdataskip6),                           //  output,    width = 1,                  .txdataskip6
		.txdataskip7              (hip_pipe_txdataskip7),                           //  output,    width = 1,                  .txdataskip7
		.rate0                    (hip_pipe_rate0),                                 //  output,    width = 2,                  .rate0
		.rate1                    (hip_pipe_rate1),                                 //  output,    width = 2,                  .rate1
		.rate2                    (hip_pipe_rate2),                                 //  output,    width = 2,                  .rate2
		.rate3                    (hip_pipe_rate3),                                 //  output,    width = 2,                  .rate3
		.rate4                    (hip_pipe_rate4),                                 //  output,    width = 2,                  .rate4
		.rate5                    (hip_pipe_rate5),                                 //  output,    width = 2,                  .rate5
		.rate6                    (hip_pipe_rate6),                                 //  output,    width = 2,                  .rate6
		.rate7                    (hip_pipe_rate7),                                 //  output,    width = 2,                  .rate7
		.rx_in0                   (hip_serial_rx_in0),                              //   input,    width = 1,        hip_serial.rx_in0
		.rx_in1                   (hip_serial_rx_in1),                              //   input,    width = 1,                  .rx_in1
		.rx_in2                   (hip_serial_rx_in2),                              //   input,    width = 1,                  .rx_in2
		.rx_in3                   (hip_serial_rx_in3),                              //   input,    width = 1,                  .rx_in3
		.rx_in4                   (hip_serial_rx_in4),                              //   input,    width = 1,                  .rx_in4
		.rx_in5                   (hip_serial_rx_in5),                              //   input,    width = 1,                  .rx_in5
		.rx_in6                   (hip_serial_rx_in6),                              //   input,    width = 1,                  .rx_in6
		.rx_in7                   (hip_serial_rx_in7),                              //   input,    width = 1,                  .rx_in7
		.tx_out0                  (hip_serial_tx_out0),                             //  output,    width = 1,                  .tx_out0
		.tx_out1                  (hip_serial_tx_out1),                             //  output,    width = 1,                  .tx_out1
		.tx_out2                  (hip_serial_tx_out2),                             //  output,    width = 1,                  .tx_out2
		.tx_out3                  (hip_serial_tx_out3),                             //  output,    width = 1,                  .tx_out3
		.tx_out4                  (hip_serial_tx_out4),                             //  output,    width = 1,                  .tx_out4
		.tx_out5                  (hip_serial_tx_out5),                             //  output,    width = 1,                  .tx_out5
		.tx_out6                  (hip_serial_tx_out6),                             //  output,    width = 1,                  .tx_out6
		.tx_out7                  (hip_serial_tx_out7),                             //  output,    width = 1,                  .tx_out7
		.npor                     (dut_npor_npor),                                  //   input,    width = 1,              npor.npor
		.pin_perst                (dut_npor_pin_perst),                             //   input,    width = 1,                  .pin_perst
		.rd_dcm_address_o         (dut_rd_dcm_master_address),                      //  output,   width = 64,     rd_dcm_master.address
		.rd_dcm_write_o           (dut_rd_dcm_master_write),                        //  output,    width = 1,                  .write
		.rd_dcm_writedata_o       (dut_rd_dcm_master_writedata),                    //  output,   width = 32,                  .writedata
		.rd_dcm_read_o            (dut_rd_dcm_master_read),                         //  output,    width = 1,                  .read
		.rd_dcm_byte_enable_o     (dut_rd_dcm_master_byteenable),                   //  output,    width = 4,                  .byteenable
		.rd_dcm_wait_request_i    (dut_rd_dcm_master_waitrequest),                  //   input,    width = 1,                  .waitrequest
		.rd_dcm_read_data_i       (dut_rd_dcm_master_readdata),                     //   input,   width = 32,                  .readdata
		.rd_dcm_read_data_valid_i (dut_rd_dcm_master_readdatavalid),                //   input,    width = 1,                  .readdatavalid
		.rd_dts_chip_select_i     (mm_interconnect_0_dut_rd_dts_slave_chipselect),  //   input,    width = 1,      rd_dts_slave.chipselect
		.rd_dts_write_i           (mm_interconnect_0_dut_rd_dts_slave_write),       //   input,    width = 1,                  .write
		.rd_dts_burst_count_i     (mm_interconnect_0_dut_rd_dts_slave_burstcount),  //   input,    width = 5,                  .burstcount
		.rd_dts_address_i         (mm_interconnect_0_dut_rd_dts_slave_address),     //   input,    width = 8,                  .address
		.rd_dts_write_data_i      (mm_interconnect_0_dut_rd_dts_slave_writedata),   //   input,  width = 256,                  .writedata
		.rd_dts_wait_request_o    (mm_interconnect_0_dut_rd_dts_slave_waitrequest), //  output,    width = 1,                  .waitrequest
		.refclk                   (refclk_clk),                                     //   input,    width = 1,            refclk.clk
		.rxm_bar2_address_o       (dut_rxm_bar2_address),                           //  output,   width = 64,          rxm_bar2.address
		.rxm_bar2_byteenable_o    (dut_rxm_bar2_byteenable),                        //  output,    width = 4,                  .byteenable
		.rxm_bar2_readdata_i      (dut_rxm_bar2_readdata),                          //   input,   width = 32,                  .readdata
		.rxm_bar2_writedata_o     (dut_rxm_bar2_writedata),                         //  output,   width = 32,                  .writedata
		.rxm_bar2_read_o          (dut_rxm_bar2_read),                              //  output,    width = 1,                  .read
		.rxm_bar2_write_o         (dut_rxm_bar2_write),                             //  output,    width = 1,                  .write
		.rxm_bar2_readdatavalid_i (dut_rxm_bar2_readdatavalid),                     //   input,    width = 1,                  .readdatavalid
		.rxm_bar2_waitrequest_i   (dut_rxm_bar2_waitrequest),                       //   input,    width = 1,                  .waitrequest
		.txs_address_i            (mm_interconnect_1_dut_txs_address),              //   input,   width = 40,               txs.address
		.txs_chipselect_i         (mm_interconnect_1_dut_txs_chipselect),           //   input,    width = 1,                  .chipselect
		.txs_byteenable_i         (mm_interconnect_1_dut_txs_byteenable),           //   input,    width = 4,                  .byteenable
		.txs_readdata_o           (mm_interconnect_1_dut_txs_readdata),             //  output,   width = 32,                  .readdata
		.txs_writedata_i          (mm_interconnect_1_dut_txs_writedata),            //   input,   width = 32,                  .writedata
		.txs_read_i               (mm_interconnect_1_dut_txs_read),                 //   input,    width = 1,                  .read
		.txs_write_i              (mm_interconnect_1_dut_txs_write),                //   input,    width = 1,                  .write
		.txs_readdatavalid_o      (mm_interconnect_1_dut_txs_readdatavalid),        //  output,    width = 1,                  .readdatavalid
		.txs_waitrequest_o        (mm_interconnect_1_dut_txs_waitrequest),          //  output,    width = 1,                  .waitrequest
		.wr_dcm_address_o         (dut_wr_dcm_master_address),                      //  output,   width = 64,     wr_dcm_master.address
		.wr_dcm_write_o           (dut_wr_dcm_master_write),                        //  output,    width = 1,                  .write
		.wr_dcm_writedata_o       (dut_wr_dcm_master_writedata),                    //  output,   width = 32,                  .writedata
		.wr_dcm_read_o            (dut_wr_dcm_master_read),                         //  output,    width = 1,                  .read
		.wr_dcm_byte_enable_o     (dut_wr_dcm_master_byteenable),                   //  output,    width = 4,                  .byteenable
		.wr_dcm_wait_request_i    (dut_wr_dcm_master_waitrequest),                  //   input,    width = 1,                  .waitrequest
		.wr_dcm_read_data_i       (dut_wr_dcm_master_readdata),                     //   input,   width = 32,                  .readdata
		.wr_dcm_read_data_valid_i (dut_wr_dcm_master_readdatavalid),                //   input,    width = 1,                  .readdatavalid
		.wr_dts_chip_select_i     (mm_interconnect_0_dut_wr_dts_slave_chipselect),  //   input,    width = 1,      wr_dts_slave.chipselect
		.wr_dts_write_i           (mm_interconnect_0_dut_wr_dts_slave_write),       //   input,    width = 1,                  .write
		.wr_dts_burst_count_i     (mm_interconnect_0_dut_wr_dts_slave_burstcount),  //   input,    width = 5,                  .burstcount
		.wr_dts_address_i         (mm_interconnect_0_dut_wr_dts_slave_address),     //   input,    width = 8,                  .address
		.wr_dts_write_data_i      (mm_interconnect_0_dut_wr_dts_slave_writedata),   //   input,  width = 256,                  .writedata
		.wr_dts_wait_request_o    (mm_interconnect_0_dut_wr_dts_slave_waitrequest)  //  output,    width = 1,                  .waitrequest
	);

	top_clk_0 clk_0 (
		.clk_out     (core_clk_out_clk),            //  output,  width = 1,          clk.clk
		.in_clk      (dut_coreclkout_hip_clk),      //   input,  width = 1,       clk_in.clk
		.reset_n     (dut_app_nreset_status_reset), //   input,  width = 1, clk_in_reset.reset_n
		.reset_n_out ()                             //  output,  width = 1,    clk_reset.reset_n
	);

	top_emif_0 emif_0 (
		.amm_ready_0         (mm_interconnect_0_emif_0_ctrl_amm_0_waitrequest),   //  output,    width = 1,       ctrl_amm_0.waitrequest_n
		.amm_read_0          (mm_interconnect_0_emif_0_ctrl_amm_0_read),          //   input,    width = 1,                 .read
		.amm_write_0         (mm_interconnect_0_emif_0_ctrl_amm_0_write),         //   input,    width = 1,                 .write
		.amm_address_0       (mm_interconnect_0_emif_0_ctrl_amm_0_address),       //   input,   width = 22,                 .address
		.amm_readdata_0      (mm_interconnect_0_emif_0_ctrl_amm_0_readdata),      //  output,  width = 512,                 .readdata
		.amm_writedata_0     (mm_interconnect_0_emif_0_ctrl_amm_0_writedata),     //   input,  width = 512,                 .writedata
		.amm_burstcount_0    (mm_interconnect_0_emif_0_ctrl_amm_0_burstcount),    //   input,    width = 7,                 .burstcount
		.amm_byteenable_0    (mm_interconnect_0_emif_0_ctrl_amm_0_byteenable),    //   input,   width = 64,                 .byteenable
		.amm_readdatavalid_0 (mm_interconnect_0_emif_0_ctrl_amm_0_readdatavalid), //  output,    width = 1,                 .readdatavalid
		.emif_usr_clk        (emif_0_emif_usr_clk_clk),                           //  output,    width = 1,     emif_usr_clk.clk
		.emif_usr_reset_n    (emif_0_emif_usr_reset_n_reset),                     //  output,    width = 1, emif_usr_reset_n.reset_n
		.global_reset_n      (dut_app_nreset_status_reset),                       //   input,    width = 1,   global_reset_n.reset_n
		.mem_ck              (emif_0_mem_mem_ck),                                 //  output,    width = 1,              mem.mem_ck
		.mem_ck_n            (emif_0_mem_mem_ck_n),                               //  output,    width = 1,                 .mem_ck_n
		.mem_a               (emif_0_mem_mem_a),                                  //  output,   width = 17,                 .mem_a
		.mem_act_n           (emif_0_mem_mem_act_n),                              //  output,    width = 1,                 .mem_act_n
		.mem_ba              (emif_0_mem_mem_ba),                                 //  output,    width = 2,                 .mem_ba
		.mem_bg              (emif_0_mem_mem_bg),                                 //  output,    width = 1,                 .mem_bg
		.mem_cke             (emif_0_mem_mem_cke),                                //  output,    width = 1,                 .mem_cke
		.mem_cs_n            (emif_0_mem_mem_cs_n),                               //  output,    width = 1,                 .mem_cs_n
		.mem_odt             (emif_0_mem_mem_odt),                                //  output,    width = 1,                 .mem_odt
		.mem_reset_n         (emif_0_mem_mem_reset_n),                            //  output,    width = 1,                 .mem_reset_n
		.mem_dqs             (emif_0_mem_mem_dqs),                                //   inout,    width = 8,                 .mem_dqs
		.mem_dqs_n           (emif_0_mem_mem_dqs_n),                              //   inout,    width = 8,                 .mem_dqs_n
		.mem_dq              (emif_0_mem_mem_dq),                                 //   inout,   width = 64,                 .mem_dq
		.mem_dbi_n           (emif_0_mem_mem_dbi_n),                              //   inout,    width = 8,                 .mem_dbi_n
		.oct_rzqin           (emif_0_oct_oct_rzqin),                              //   input,    width = 1,              oct.oct_rzqin
		.pll_ref_clk         (emif_0_pll_ref_clk_clk),                            //   input,    width = 1,      pll_ref_clk.clk
		.local_cal_success   (emif_0_status_local_cal_success),                   //  output,    width = 1,           status.local_cal_success
		.local_cal_fail      (emif_0_status_local_cal_fail)                       //  output,    width = 1,                 .local_cal_fail
	);

	top_onchip_memory2_0 onchip_memory2_0 (
		.clk         (dut_coreclkout_hip_clk),                           //   input,    width = 1,   clk1.clk
		.clk2        (dut_coreclkout_hip_clk),                           //   input,    width = 1,   clk2.clk
		.reset       (rst_controller_reset_out_reset),                   //   input,    width = 1, reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),               //   input,    width = 1,       .reset_req
		.reset2      (rst_controller_reset_out_reset),                   //   input,    width = 1, reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req),               //   input,    width = 1,       .reset_req
		.address     (mm_interconnect_0_onchip_memory2_0_s1_address),    //   input,   width = 11,     s1.address
		.clken       (mm_interconnect_0_onchip_memory2_0_s1_clken),      //   input,    width = 1,       .clken
		.chipselect  (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //   input,    width = 1,       .chipselect
		.write       (mm_interconnect_0_onchip_memory2_0_s1_write),      //   input,    width = 1,       .write
		.readdata    (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //  output,  width = 256,       .readdata
		.writedata   (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //   input,  width = 256,       .writedata
		.byteenable  (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //   input,   width = 32,       .byteenable
		.address2    (mm_interconnect_0_onchip_memory2_0_s2_address),    //   input,   width = 11,     s2.address
		.chipselect2 (mm_interconnect_0_onchip_memory2_0_s2_chipselect), //   input,    width = 1,       .chipselect
		.clken2      (mm_interconnect_0_onchip_memory2_0_s2_clken),      //   input,    width = 1,       .clken
		.write2      (mm_interconnect_0_onchip_memory2_0_s2_write),      //   input,    width = 1,       .write
		.readdata2   (mm_interconnect_0_onchip_memory2_0_s2_readdata),   //  output,  width = 256,       .readdata
		.writedata2  (mm_interconnect_0_onchip_memory2_0_s2_writedata),  //   input,  width = 256,       .writedata
		.byteenable2 (mm_interconnect_0_onchip_memory2_0_s2_byteenable)  //   input,   width = 32,       .byteenable
	);

	top_hw_altera_mm_interconnect_191_scrfrry mm_interconnect_0 (
		.DUT_dma_rd_master_address                                      (dut_dma_rd_master_address),                         //   input,   width = 64,                                        DUT_dma_rd_master.address
		.DUT_dma_rd_master_waitrequest                                  (dut_dma_rd_master_waitrequest),                     //  output,    width = 1,                                                         .waitrequest
		.DUT_dma_rd_master_burstcount                                   (dut_dma_rd_master_burstcount),                      //   input,    width = 5,                                                         .burstcount
		.DUT_dma_rd_master_byteenable                                   (dut_dma_rd_master_byteenable),                      //   input,   width = 32,                                                         .byteenable
		.DUT_dma_rd_master_write                                        (dut_dma_rd_master_write),                           //   input,    width = 1,                                                         .write
		.DUT_dma_rd_master_writedata                                    (dut_dma_rd_master_writedata),                       //   input,  width = 256,                                                         .writedata
		.DUT_dma_wr_master_address                                      (dut_dma_wr_master_address),                         //   input,   width = 64,                                        DUT_dma_wr_master.address
		.DUT_dma_wr_master_waitrequest                                  (dut_dma_wr_master_waitrequest),                     //  output,    width = 1,                                                         .waitrequest
		.DUT_dma_wr_master_burstcount                                   (dut_dma_wr_master_burstcount),                      //   input,    width = 5,                                                         .burstcount
		.DUT_dma_wr_master_read                                         (dut_dma_wr_master_read),                            //   input,    width = 1,                                                         .read
		.DUT_dma_wr_master_readdata                                     (dut_dma_wr_master_readdata),                        //  output,  width = 256,                                                         .readdata
		.DUT_dma_wr_master_readdatavalid                                (dut_dma_wr_master_readdatavalid),                   //  output,    width = 1,                                                         .readdatavalid
		.DUT_rxm_bar2_address                                           (dut_rxm_bar2_address),                              //   input,   width = 64,                                             DUT_rxm_bar2.address
		.DUT_rxm_bar2_waitrequest                                       (dut_rxm_bar2_waitrequest),                          //  output,    width = 1,                                                         .waitrequest
		.DUT_rxm_bar2_byteenable                                        (dut_rxm_bar2_byteenable),                           //   input,    width = 4,                                                         .byteenable
		.DUT_rxm_bar2_read                                              (dut_rxm_bar2_read),                                 //   input,    width = 1,                                                         .read
		.DUT_rxm_bar2_readdata                                          (dut_rxm_bar2_readdata),                             //  output,   width = 32,                                                         .readdata
		.DUT_rxm_bar2_readdatavalid                                     (dut_rxm_bar2_readdatavalid),                        //  output,    width = 1,                                                         .readdatavalid
		.DUT_rxm_bar2_write                                             (dut_rxm_bar2_write),                                //   input,    width = 1,                                                         .write
		.DUT_rxm_bar2_writedata                                         (dut_rxm_bar2_writedata),                            //   input,   width = 32,                                                         .writedata
		.emif_0_ctrl_amm_0_address                                      (mm_interconnect_0_emif_0_ctrl_amm_0_address),       //  output,   width = 22,                                        emif_0_ctrl_amm_0.address
		.emif_0_ctrl_amm_0_write                                        (mm_interconnect_0_emif_0_ctrl_amm_0_write),         //  output,    width = 1,                                                         .write
		.emif_0_ctrl_amm_0_read                                         (mm_interconnect_0_emif_0_ctrl_amm_0_read),          //  output,    width = 1,                                                         .read
		.emif_0_ctrl_amm_0_readdata                                     (mm_interconnect_0_emif_0_ctrl_amm_0_readdata),      //   input,  width = 512,                                                         .readdata
		.emif_0_ctrl_amm_0_writedata                                    (mm_interconnect_0_emif_0_ctrl_amm_0_writedata),     //  output,  width = 512,                                                         .writedata
		.emif_0_ctrl_amm_0_burstcount                                   (mm_interconnect_0_emif_0_ctrl_amm_0_burstcount),    //  output,    width = 7,                                                         .burstcount
		.emif_0_ctrl_amm_0_byteenable                                   (mm_interconnect_0_emif_0_ctrl_amm_0_byteenable),    //  output,   width = 64,                                                         .byteenable
		.emif_0_ctrl_amm_0_readdatavalid                                (mm_interconnect_0_emif_0_ctrl_amm_0_readdatavalid), //   input,    width = 1,                                                         .readdatavalid
		.emif_0_ctrl_amm_0_waitrequest                                  (~mm_interconnect_0_emif_0_ctrl_amm_0_waitrequest),  //   input,    width = 1,                                                         .waitrequest
		.DUT_rd_dts_slave_address                                       (mm_interconnect_0_dut_rd_dts_slave_address),        //  output,    width = 8,                                         DUT_rd_dts_slave.address
		.DUT_rd_dts_slave_write                                         (mm_interconnect_0_dut_rd_dts_slave_write),          //  output,    width = 1,                                                         .write
		.DUT_rd_dts_slave_writedata                                     (mm_interconnect_0_dut_rd_dts_slave_writedata),      //  output,  width = 256,                                                         .writedata
		.DUT_rd_dts_slave_burstcount                                    (mm_interconnect_0_dut_rd_dts_slave_burstcount),     //  output,    width = 5,                                                         .burstcount
		.DUT_rd_dts_slave_waitrequest                                   (mm_interconnect_0_dut_rd_dts_slave_waitrequest),    //   input,    width = 1,                                                         .waitrequest
		.DUT_rd_dts_slave_chipselect                                    (mm_interconnect_0_dut_rd_dts_slave_chipselect),     //  output,    width = 1,                                                         .chipselect
		.onchip_memory2_0_s2_address                                    (mm_interconnect_0_onchip_memory2_0_s2_address),     //  output,   width = 11,                                      onchip_memory2_0_s2.address
		.onchip_memory2_0_s2_write                                      (mm_interconnect_0_onchip_memory2_0_s2_write),       //  output,    width = 1,                                                         .write
		.onchip_memory2_0_s2_readdata                                   (mm_interconnect_0_onchip_memory2_0_s2_readdata),    //   input,  width = 256,                                                         .readdata
		.onchip_memory2_0_s2_writedata                                  (mm_interconnect_0_onchip_memory2_0_s2_writedata),   //  output,  width = 256,                                                         .writedata
		.onchip_memory2_0_s2_byteenable                                 (mm_interconnect_0_onchip_memory2_0_s2_byteenable),  //  output,   width = 32,                                                         .byteenable
		.onchip_memory2_0_s2_chipselect                                 (mm_interconnect_0_onchip_memory2_0_s2_chipselect),  //  output,    width = 1,                                                         .chipselect
		.onchip_memory2_0_s2_clken                                      (mm_interconnect_0_onchip_memory2_0_s2_clken),       //  output,    width = 1,                                                         .clken
		.DUT_wr_dts_slave_address                                       (mm_interconnect_0_dut_wr_dts_slave_address),        //  output,    width = 8,                                         DUT_wr_dts_slave.address
		.DUT_wr_dts_slave_write                                         (mm_interconnect_0_dut_wr_dts_slave_write),          //  output,    width = 1,                                                         .write
		.DUT_wr_dts_slave_writedata                                     (mm_interconnect_0_dut_wr_dts_slave_writedata),      //  output,  width = 256,                                                         .writedata
		.DUT_wr_dts_slave_burstcount                                    (mm_interconnect_0_dut_wr_dts_slave_burstcount),     //  output,    width = 5,                                                         .burstcount
		.DUT_wr_dts_slave_waitrequest                                   (mm_interconnect_0_dut_wr_dts_slave_waitrequest),    //   input,    width = 1,                                                         .waitrequest
		.DUT_wr_dts_slave_chipselect                                    (mm_interconnect_0_dut_wr_dts_slave_chipselect),     //  output,    width = 1,                                                         .chipselect
		.onchip_memory2_0_s1_address                                    (mm_interconnect_0_onchip_memory2_0_s1_address),     //  output,   width = 11,                                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                      (mm_interconnect_0_onchip_memory2_0_s1_write),       //  output,    width = 1,                                                         .write
		.onchip_memory2_0_s1_readdata                                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),    //   input,  width = 256,                                                         .readdata
		.onchip_memory2_0_s1_writedata                                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),   //  output,  width = 256,                                                         .writedata
		.onchip_memory2_0_s1_byteenable                                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),  //  output,   width = 32,                                                         .byteenable
		.onchip_memory2_0_s1_chipselect                                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),  //  output,    width = 1,                                                         .chipselect
		.onchip_memory2_0_s1_clken                                      (mm_interconnect_0_onchip_memory2_0_s1_clken),       //  output,    width = 1,                                                         .clken
		.onchip_memory2_0_reset2_reset_bridge_in_reset_reset            (rst_controller_reset_out_reset),                    //   input,    width = 1,            onchip_memory2_0_reset2_reset_bridge_in_reset.reset
		.emif_0_ctrl_amm_0_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                //   input,    width = 1, emif_0_ctrl_amm_0_translator_reset_reset_bridge_in_reset.reset
		.DUT_coreclkout_hip_clk                                         (dut_coreclkout_hip_clk),                            //   input,    width = 1,                                       DUT_coreclkout_hip.clk
		.emif_0_emif_usr_clk_clk                                        (emif_0_emif_usr_clk_clk)                            //   input,    width = 1,                                      emif_0_emif_usr_clk.clk
	);

	top_hw_altera_mm_interconnect_191_3pabmzq mm_interconnect_1 (
		.DUT_rd_dcm_master_address                                      (dut_rd_dcm_master_address),               //   input,  width = 64,                                        DUT_rd_dcm_master.address
		.DUT_rd_dcm_master_waitrequest                                  (dut_rd_dcm_master_waitrequest),           //  output,   width = 1,                                                         .waitrequest
		.DUT_rd_dcm_master_byteenable                                   (dut_rd_dcm_master_byteenable),            //   input,   width = 4,                                                         .byteenable
		.DUT_rd_dcm_master_read                                         (dut_rd_dcm_master_read),                  //   input,   width = 1,                                                         .read
		.DUT_rd_dcm_master_readdata                                     (dut_rd_dcm_master_readdata),              //  output,  width = 32,                                                         .readdata
		.DUT_rd_dcm_master_readdatavalid                                (dut_rd_dcm_master_readdatavalid),         //  output,   width = 1,                                                         .readdatavalid
		.DUT_rd_dcm_master_write                                        (dut_rd_dcm_master_write),                 //   input,   width = 1,                                                         .write
		.DUT_rd_dcm_master_writedata                                    (dut_rd_dcm_master_writedata),             //   input,  width = 32,                                                         .writedata
		.DUT_wr_dcm_master_address                                      (dut_wr_dcm_master_address),               //   input,  width = 64,                                        DUT_wr_dcm_master.address
		.DUT_wr_dcm_master_waitrequest                                  (dut_wr_dcm_master_waitrequest),           //  output,   width = 1,                                                         .waitrequest
		.DUT_wr_dcm_master_byteenable                                   (dut_wr_dcm_master_byteenable),            //   input,   width = 4,                                                         .byteenable
		.DUT_wr_dcm_master_read                                         (dut_wr_dcm_master_read),                  //   input,   width = 1,                                                         .read
		.DUT_wr_dcm_master_readdata                                     (dut_wr_dcm_master_readdata),              //  output,  width = 32,                                                         .readdata
		.DUT_wr_dcm_master_readdatavalid                                (dut_wr_dcm_master_readdatavalid),         //  output,   width = 1,                                                         .readdatavalid
		.DUT_wr_dcm_master_write                                        (dut_wr_dcm_master_write),                 //   input,   width = 1,                                                         .write
		.DUT_wr_dcm_master_writedata                                    (dut_wr_dcm_master_writedata),             //   input,  width = 32,                                                         .writedata
		.DUT_txs_address                                                (mm_interconnect_1_dut_txs_address),       //  output,  width = 40,                                                  DUT_txs.address
		.DUT_txs_write                                                  (mm_interconnect_1_dut_txs_write),         //  output,   width = 1,                                                         .write
		.DUT_txs_read                                                   (mm_interconnect_1_dut_txs_read),          //  output,   width = 1,                                                         .read
		.DUT_txs_readdata                                               (mm_interconnect_1_dut_txs_readdata),      //   input,  width = 32,                                                         .readdata
		.DUT_txs_writedata                                              (mm_interconnect_1_dut_txs_writedata),     //  output,  width = 32,                                                         .writedata
		.DUT_txs_byteenable                                             (mm_interconnect_1_dut_txs_byteenable),    //  output,   width = 4,                                                         .byteenable
		.DUT_txs_readdatavalid                                          (mm_interconnect_1_dut_txs_readdatavalid), //   input,   width = 1,                                                         .readdatavalid
		.DUT_txs_waitrequest                                            (mm_interconnect_1_dut_txs_waitrequest),   //   input,   width = 1,                                                         .waitrequest
		.DUT_txs_chipselect                                             (mm_interconnect_1_dut_txs_chipselect),    //  output,   width = 1,                                                         .chipselect
		.DUT_rd_dcm_master_translator_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),          //   input,   width = 1, DUT_rd_dcm_master_translator_reset_reset_bridge_in_reset.reset
		.DUT_coreclkout_hip_clk                                         (dut_coreclkout_hip_clk)                   //   input,   width = 1,                                       DUT_coreclkout_hip.clk
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~dut_app_nreset_status_reset),       //   input,  width = 1, reset_in0.reset
		.clk            (dut_coreclkout_hip_clk),             //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     //  output,  width = 1, reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //  output,  width = 1,          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~emif_0_emif_usr_reset_n_reset),     //   input,  width = 1, reset_in0.reset
		.clk            (emif_0_emif_usr_clk_clk),            //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

endmodule
